library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use IEEE.std_logic_textio.all;          -- I/O for logic types
library STD;
use STD.textio.all;                     -- basic I/O
use work.types.all;
 
entity convolution_engine_tb is
end convolution_engine_tb;
 
architecture behavior of convolution_engine_tb is
    -- Component Declaration for the Unit Under Test (UUT)
    component convolution_engine
        port(
            clk         : in  STD_LOGIC;
            rst         : in  STD_LOGIC;
            new_data    : in  STD_LOGIC;          
            data_input  : in  STD_LOGIC_VECTOR(AXIS_BUS_WIDTH - 1 downto 0);
            done        : out STD_LOGIC;         
            conv_output : out STD_LOGIC_VECTOR(AXIS_BUS_WIDTH - 1 downto 0)
        );
    end component;

    -- Inputs
    signal clk        : std_logic := '0';
    signal rst        : std_logic := '0';
    signal new_data   : std_logic := '0';
    signal data_input : std_logic_vector(AXIS_BUS_WIDTH - 1 downto 0) := (others => '0');

    -- Outputs
    signal done        : STD_LOGIC := '0';
    signal conv_output : STD_LOGIC_VECTOR(AXIS_BUS_WIDTH - 1 downto 0) := (others => '0');
--    signal conv_output : tp_act_value_mem_data := (others => (others => '0'));

    -- Clock period definitions
    constant clk_period : time := 1 ns;
begin
    -- Instantiate the Unit Under Test (UUT)
    uut: convolution_engine
        port map(
            clk => clk,
            rst => rst,
            new_data => new_data,
            data_input => data_input,
            done => done,
            conv_output => conv_output
        );

    -- Clock process definitions
    clk_process: process
    begin
        clk <= '1';
        wait for clk_period/2;

        clk <= '0';
        wait for clk_period/2;
    end process;

    -- Stimulus process
    stim_proc: process
        variable my_line : line;  -- type 'line' comes from textio
    begin
        -- hold reset state for 10 ns.
        rst <= '1';
        wait for 10 ns;

        rst <= '0';

        ---------------------------------------
        -- Image to process from DDR to BRAM --
        ---------------------------------------
        -- Indices #transfers - 1
        new_data <= '1';
        data_input <= "00000000000000000000101111010000";
        wait for clk_period;

        -- Indices
        new_data <= '1';
        data_input <= "11111011111111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011111110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011111101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10111011111101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011111110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11011011111111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011110111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11001011110111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10001011111111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11011011111110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011111110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011111111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011111111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011111111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011111110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011111110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101011111110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10101011101111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11011011111110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011111110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10011011111110010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11011011111110010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10101011101111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011111110010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101111101110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10001011111111010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11001011111110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10001011111111010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11001011111110010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10001011101111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10111011111111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011111110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10101011111111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00111011111111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111101111110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11001101101110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10101011101111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10111011111111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111001111110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101011111111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10111011111111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011111110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10101011111101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101011111101010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101011111100010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101011111101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10101011111101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10101011111101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011111110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011111110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101011111100110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101111111100110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111111111100110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111111111101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10101111111101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10111011111101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011111101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011111110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011111111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10111011111111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011111110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011111111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10101011110111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011111110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011111110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011111110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10111011111111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011111110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011111110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011111110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10111011110111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11011011110110010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101011101111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10011011111111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11011011111110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10001011111110010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11001011111110010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10001111101111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101011111110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101111101110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10001011111111010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11001011111110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10001011111111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11001011111110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10101011101111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10111011111111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111001111110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10101011111111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "01111011111111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111001111110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101101101110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10001011111111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011111111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011111110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10101011111111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011111110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10111011111101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10101011111101010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101011111100010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101011111100110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10101011111101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00101011111111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011111110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011111110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101111111100110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101111111100110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101011111101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10101111111101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10101111111101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10111111111111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101011110100110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10101011101101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10111011111101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10111011111101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011111110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011111111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011111111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011111111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11001011110110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11001011110110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011111110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10111011111111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101011111111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011111110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011111110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10101011111111010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11011011110110010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11001011111110010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10101011111111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011111110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011111110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11001011111110010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101011101111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011111111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101111111110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10001011101111010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11001011111110010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10001011101111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11001011111111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10101011101111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10111011111111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011111110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10001011111111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "01111011111110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111001111110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101111101110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10001011111111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011111110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011101111010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10101011111111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011111110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10101011111101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10101011111100010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101011111110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10101011111111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10101011111101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011111111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111111111110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101111111110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101011111100110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10101011111101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10101111111101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10111111111101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10111111111111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111111111111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011111100110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011111100110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101011101111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10001011111101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101011111100110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11011011111110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10111011111111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011111110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10011011111111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11001011110110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11001011110110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10011011110111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10001011110111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011111110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011110110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10001011101111010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10001011110111010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11011011111110010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10101011101111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101011111110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011111110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101011111110010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11001011101110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10001011111111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11001111111110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10101011101111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11001011111110010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11001011101111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10001011111111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101011101111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10111011111111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011111110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10101011111111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011111110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111001101110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11001011101110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10001011111111010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011111110010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10001011111111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00111011111111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011111110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10101011111101010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101011111100010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10101011111111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10101011111101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10101011111101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111111111100110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101101111100110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101111111100110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10101111111101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10101011111101010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10111011111101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111111111101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111111111101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111111111111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011111100110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011111100110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011111110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101011111111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10001011101111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11011011111110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11011011101110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10101011111111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011111111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11011011110110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11001011110110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11011011110111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10011011110111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10101011110110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011110110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011111110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10101011111111010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101011111110010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101011111110010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10101011111111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011111110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101011101110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101111101110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10001111111111010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11001111111110010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101011101110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11001111101110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10001011101111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10001011111111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10101011101111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10001011111110010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101011101110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10101011111111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011111110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101011101110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10001011111110010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10001011101111010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101011111110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10101011111111010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10111011111111010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011111101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101011111100010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101011111100110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10101011111101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10101011111101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111111111100110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101001111100110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101011101100110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10101111111101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10101011111101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00111111111101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10111111111101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111111111110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111111111110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011111101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011111101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011111101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011111110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011111110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011111110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10101011101111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11001011101110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10101011101111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10011011111111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11011011110111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011110110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11011011110110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11011011110110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10001011110111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11011011110110010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11011011110110010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101111101111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101111111111010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101011111111010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10101011111111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11011011111110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101011111110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101111101110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10101011101111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101111111110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11001011101110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10001011111111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11001011101110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10001111101111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10001011101111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11001011111110010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101011101110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10101011111111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011111110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10101011101111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11001011111110010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11001011101110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101011101110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10001011101111010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101011111110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101011111101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011111100110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10101011111101010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10101011111101010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101011111100110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011111100010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101011101100010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101111111101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10101111111101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00111011111101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111111111101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111111111111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111111111101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111111111100110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101011111100110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011111111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111111111111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011111111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011111110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011111110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101011111110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10101011101111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101011111101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10101011111111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10101011110111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10011011110110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11011011110110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11011011110110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11011011110111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10101011110111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101011110110010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101011111110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101111111111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101111101110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10101011101111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101011111111010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101011111110010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101011101110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10101011101111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11001011111111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11001011101110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10001011101111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11001011101110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10001111101111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10101111101111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101111101110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10101011101111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10111011111111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011111110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10001011111111010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11001011111110010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101011101110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101111101110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10101011101111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10101011111111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101011111100010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011111110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10101011111101010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10101011111101010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011111100110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101011111100110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101111111101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10101111111101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10111111111101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10111011111111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111111111110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111111111100110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101111111100110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111111111100110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111111111101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10111011111101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10111011111101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011111101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011111111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011111110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101011111110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10101011111111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10101011111101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011111111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011111110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10001011110111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11011011110110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101011111111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011111110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101011101111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101011111101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011111100110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101011101111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101011111111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101011101111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10101011111111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101011111110010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101011101110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11001011101110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10101111111111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11001011111110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10101011101111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11001011111110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101111101111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10101011101111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101011111110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10101011101111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10001011111111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111111111110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10001011111111010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11001011111110010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101011101110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101111101110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10101011111111010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011111101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011111110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101011101110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10101011111101010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011111100110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011111100110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101011111101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00101111111101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00111111111101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111111111101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111111111100110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111111111100110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111111111100110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111111111100110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10101111111101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10111111111101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011111101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10101011111101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10101011111101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10111011111111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "01111011111111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011111110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101011111110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10101011111111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011111110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011111110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10101011101111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10101011111111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00101011111101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "01111011111110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011111110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10101011111101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "01111011111100110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011111110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101011101111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101111101110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10101011101111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11001011111110010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11001011101111010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11001011101110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10101011101111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101011111110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101011101111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11001011111110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101011101111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11001011101110010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101111101110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101011101111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10001011111111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101111111110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10001011101110010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11001011101110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101011101110010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11001011101111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10101011111111010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011111110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011111110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10101111111111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011111100010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011111100110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011111101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00101011111101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00111111111111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111111111111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111101111100110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111111111100110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101111111100110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101111111101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011111101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10111011111101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10111111111101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "01111011111100110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011111100110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011111101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10101011111101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10111011111101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011111101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011111110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011111110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011111110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10101011111101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "01111011111101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011111110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10111011111111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011111100110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011111110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10111011111111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011111111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011111110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101011101111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101011111110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10101011101111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101011111111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101011101110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10101011101110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10101011101111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101011111110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101011101111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11001011111110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10101011101111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11001011101110010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10101111101111010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10101111101111010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10001011111111010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101011111110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101011101110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10101011101111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "01101011111110010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101011101111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10111011111111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011111110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011111111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101011111101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011111100110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011111101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10101011111101010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00111111111111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111111111110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111101111100110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111111111100110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111111111110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10101111111111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10111011111101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011111101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011111101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101011111101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111111111110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "01111011111100110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011111110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011111111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10111011101101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10111011111111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011111111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011111110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011111100110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101011111101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011111101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111001101110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101111101110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101111101111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101011111110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101011101110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10101111101111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011101110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101011101111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101011111111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101011101111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101011111111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101011111110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10001011101110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10001011101110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11001011101110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11001011101111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11001011101110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10101011101111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11001011101110010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10101011101111010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10001111101111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10001011111111010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11001011111110010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11001011101110010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10101011111111010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101011111110010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10101011111111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011111111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011111111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10101011111111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011111111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011111101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10101011111101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00101011111101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111111111100110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111101111100110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111111111100110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011111101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111111111101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111111111100110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101011111100110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111111111101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101111111101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111111111101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10111011111101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011111101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011111110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "01111011111110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011111110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011111111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10101011101101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10101011111101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011111110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101011111110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101011101110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101011101111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101111101110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101111101111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10101111101111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101111101111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101111101111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101111101111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101111101111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101011101111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101011101110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101011101111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101011111111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11001011101110010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10001011101110010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10001011101110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10001011101111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11001011111110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10001011101111010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11001011101110010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11001111101110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10001111101111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101011111111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11001111101110010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10001011101110010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10101011111111010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101011101110010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10101011111111010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011111110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10101011111111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101011111111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011111100110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10101011111101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00101011111101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111111111100110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111101111100110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011111100110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101111111101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111111111100110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101111111101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101111111101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101111111101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "01101111111101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00101111111101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "01111111111101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011111101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101011111111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10101011111111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10111011110111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011111110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011111110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011111111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10111011101111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10111011111101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11011011111100110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11001011110110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101011111110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10101011101111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101111101110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101011101111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101111101111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101111101110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10101111101111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101011101111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101011101111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101011101110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101011101111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101011101111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11001011101110010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10001011111111010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11001011101110010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10101011101111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011111110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11011011111110010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11001011111110010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11011011101110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10001111101111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101011111111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11001011101110010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10001011101110010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101011101110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10101011101111010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10111011111101010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101011101111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10111011111111010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011111110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101011111101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10101011111101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011111101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111101111100110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111101101100110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101111101100110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101111111101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101111111101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00101111111101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "01101111111101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "01111111111101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111111111111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111111111111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111111111111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011111100110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011111100110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011111101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10101011111101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10101011111101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011111101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011111110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011111110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011111111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10001011110101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11011011111100110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101111111110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101111101111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101011101111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101111101110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101111101111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101011101111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101111101111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101011101111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101011101110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101011101110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11001011101110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10001011111111010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11001011111110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10001011111111010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11011011111110010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10111011111111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "01111011111110010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11011011111110010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011111110010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011101110010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10001111111111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11011011111110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11001011101110010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101011101110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101111101110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10101011101111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101011101111010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10101011101111010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101011111101010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101011101111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10101011111101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011111101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111101111100110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111101101100110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101111111101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10101111111101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00101111111101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "01111111111101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111111111111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111111111100110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011111100110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111111111111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101111111111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111111111101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011111111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011111101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011111100110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011111110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011101111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10101111101111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10101011111101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011111101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11011011110100110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11001011111110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10001011101111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11001111111111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101011111110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101011111110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101011101111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101111101110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101011101111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11001011100110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101111101111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101111101110010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101011101110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10101011101101010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10101011111111010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101011111110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10001011111111010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011111110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10111011101111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011111110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11011011101110010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011101110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011101111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10111011111111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011111110010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11011011111110010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011101110010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101111101110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101111101111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101111101111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10101011111111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101011101111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10101011111111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10111011111101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111101111100110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111101101110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10101011111111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10101111111101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00111111111101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111111111101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111101111100110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101101111100110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101101101100110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101111101101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10101111111101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10101011111101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101111111101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101011101101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101011101101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10111011111101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011111101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011111100110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011111111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011101111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10101011111111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011111100110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11011011110100110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11001011111110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10001111101111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101011111110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101011111110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101011101111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101011101111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101011101110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11001011100110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101011101110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10101011101111010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10101011101110010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10001111111111010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011111110010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10111011101110010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11001011101110010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11001011101110010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10001011101111010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11011111101110010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111111101110010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011101110010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10111011101111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10111011111111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11011011111110010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011111100010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011111110010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111111101110010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101111101110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10101111101101010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101011101101010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10101011101101010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10101011111101010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011111100110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111111101100110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10101011111101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00101011111101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011111101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111101111100110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111101111100110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101101101100110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101101101110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101111101111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10101111101101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10101111111101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101111111101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10101111111101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "01111011111100110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101011111100110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101011101101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10101011111101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10111011111101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011111101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011111100110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011111110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101111101111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101011111111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101011111110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101111101111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101111101111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101011110111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101111111110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101011101111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101011101111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101111101110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101111100110010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10101011101111010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10101011101111010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10001111101110010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11001011101110010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011101110010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11001011101110010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10001011101110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10001011101111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11011011101110010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10111011101111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011101110010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10011011101111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10011011101111010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011101100010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10111011111101010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011111010010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011101100010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111111101110010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101111101111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101111101111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10101011101101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10101011111101010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101111101100110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10101011111101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10111011111101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101011111101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111101111100110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101101101100110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101111101110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101111101101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101111111101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "01101111111101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "01101111111101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "01101011111101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "01101111111101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101111111101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011111101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011110101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "01111011111100110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101011111100110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101011101111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10101011111101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10111011111101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011111101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011111100110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011111111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10101011101111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101011111101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101011101100110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101011100101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101011100111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101111101110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101011101111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10101111101101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101111111111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011111110010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011101110010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10001011101110010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11001011101110010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11011011101110010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101011101110010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10011111101110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10111011101111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11011011101110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10011011101111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11011011101110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10111111101111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011101111010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111111101111010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10101011101101010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011111100010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111111111100010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111111101100110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111111101100010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10101111101101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101011101101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101111101100110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10101111111101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10101111111101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101111111101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101101101100110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101111101110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101111101111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10101111111101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00101111111101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "01101111111101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101111111101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111111111100110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111111111100110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111111111101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111111111101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10101011100101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10101011110101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011111101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011111100110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011111100110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011111110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10101011101111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10111011111111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011111111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011111100110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011111100110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101011100101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101011111101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101011101100110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101011100111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101011101111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101011111100110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10101111101111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10101011111111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011111110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011101110010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10111011101111010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10011011101111010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11011011101110010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11011111101110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10011111101111010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10011111101111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11011111101110010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11011011101110010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011101110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10111111101111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011101110010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10101111101111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101111101101010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10111011101101010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10111011111111010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111111111100010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111111101100110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101111101101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101111101100110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10101111101101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10101111111101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101111111101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101111101110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101111101111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00101111111101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "01101111111101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101111111101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101111111100110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101111111100110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101111101100110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111111101101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101111111101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00111111111101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00111111111101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101111100101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101111101101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10101011101101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10101011101101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10111011111101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011111100110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011111110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011101111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10101011101111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011111100110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011111100110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101011111110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101111101111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101111101100110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101111101101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101011101101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10101011101101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10101011111111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011111110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011101110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011101110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111111101110010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10011011101111010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11011011101110010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11011111101110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10011111101111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11011111101110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10011111101111010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011101110010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111111101110010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10111111101111010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10111111101111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10111111101111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10111111101101010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10111011101101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10111011111111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111111111010110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111111101100010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111111101100010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10101111101101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10101111111101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101111101101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101111101110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10101111111101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10101111111101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101111111101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101111111100110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101111101100110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101111111101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "01101111111101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "01101111111101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "01111111111101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00111111111101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00111111111101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111111111111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "01111011111100110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "01111011111100110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101011111101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101111111111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101011101111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10101011101111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10111011111111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011111111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011111110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011111101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011111111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101011111100110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101011111100110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101111101101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101111111111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101111111111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101011101111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10101011101111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10111011101111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011101110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011101110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11011111101110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11011111101111010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111111101110010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11011111101110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10011111101111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11011111101110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10011111101111010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011101110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111111101110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10011111101111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10111011101111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111111101110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10111111101101010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10101111101101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10111011101111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011111100110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111111101100010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111111101101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101111101101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101111101101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101111101110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101111101101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10101111111101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101111111101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101111101100110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101111111101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10101111111101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00101111111101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00111111111101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111111111101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111111111101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111111111101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111111111101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111111111101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011111101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011111101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101011111101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101011111100110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101111111100110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101011111110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10101011101111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10101011101111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10111011111101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011111101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011111110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011101111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101011101101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101111101100110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101111101101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10101011101111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101011111101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011111100110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011100110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10111011101111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011101110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11011111101110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111111101111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10011111101111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11011111101110010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10011111101111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11011111101110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10011111101111010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111111101110010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11011111101110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10111111101111010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10111011101111010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111111101100110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10101111101101010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111111101101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111111101100110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111111101101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111111111101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111111111101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111111101100110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101111101100110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101111101111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10101111101101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101111101101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101111101101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00101111111101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00101111111101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111111111101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111111111101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111111111100110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101101111100110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101111101101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101111111101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101111101101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101111111101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101011101101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101011101101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101011101101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10111011110101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011110101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "01111011111101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011111100110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111111111111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10011011101101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10111011111101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011111100110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011111100110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101111111100110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101011101101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10101011101101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10101011100111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10101011111111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011111110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011100110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011101110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10111011101111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111111100110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111111101110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10011111101111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11011111101110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10011011101111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11011111101110010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10111111101111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111111101110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111111101111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10111111101111010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10111011101111010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111111101110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10111111101101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111101101100010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111111101101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10111011101111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00111011111101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111111111100110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111111101100110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101111101101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101111101111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101111101111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101111101111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10101111101101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10101111111101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101111111101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101101111100110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101101101100110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101111101101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101111101101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101111111101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "01101111111101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "01101111111101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "01101111111101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101111111111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101111101111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101011101101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10101011100101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10101011110101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10111011111101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011111101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011111101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011111100110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111111101111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10111011101111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011111100110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101011111100110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101111101100110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101011101101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10101011101101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10111011111101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011101100110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011101110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011100110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011101110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011101111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111111101110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111111101111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111111101111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10111111101111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11011111101110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111111101111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111111101110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111111101111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10111111101111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10111011101111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111111101110010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10111111101100010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111111101101010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10111111101101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10101111101111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011111111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111111111100110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111111111100110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101111101101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101111101111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10101111111101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "01101111111101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101111101101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101111101101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101111101101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101111111101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10101111111101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00101111111101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "01101111111101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "01101111111101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "01101111111101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011111101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011111101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "01111011111101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011111101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "01101011111101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "01101011111101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101111101111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10101011101111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10101011101101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10111011111101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011111101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011111100110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111111111100110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111111111100110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111111101101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101011101100110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101011100101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011100101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011100101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011100100110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111111101111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10111011101111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011101100110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011100100110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111111100110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111111101110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10111111101111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111111101111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111111101110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111111101111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111111101111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111111101111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10111111101111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10111111101111010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111111101101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111111101101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111111101101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10111111101101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10111111101101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10111111101101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011111100110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111111101100110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101111101111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10101111111101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101111111101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101111111100110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101111101100110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10101111111101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00101111111101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00101111111101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10111111111101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011111101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111111111101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011111101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011111101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011111101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011111101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101011100101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101011100101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10101011111101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011111101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101011111101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101011111100110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101111111111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101011101111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10101011101101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10111011111101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011111100110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011111100110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011111100110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101111101101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101011100101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011110100110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011110100110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011100100110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111111101101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111111101101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111111101101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111111101100110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111111101110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111111101110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10111111101111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10111111101111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111111101110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10111111101111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011101110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111111101110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10111111101111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10111111101111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111111101110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10111111101111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111111101101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111111101101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111111101101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10111011101101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111111101100110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111111101101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111111101101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101111101101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101111101101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101111101101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101111111101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101111110101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101011111101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101011111101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101111111101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101101111101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101101101101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101101101101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10101111101101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101011111101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101011111101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101111101101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101111101111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101111101111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10101011101111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10101011101101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101011101101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10101011101101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10101011111101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011111100110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011111100110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111111101111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111111101111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111111101100110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101111100100110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101111101101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011100101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011100100110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111111100101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111111101101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111111100101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11011111100111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11011111101111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111111101110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111111101111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111111101111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10111111101111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111111101110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10111011101111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011111110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011101110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111111101111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111111101111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10111111101111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10111111101101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10111111101101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111111101111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111111101111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10111011101101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011101100110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111111101101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10101111111101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00101111111101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "01101111111101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "01101111111101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101111111101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101111101100110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101111101101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101111101111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101111101101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101111101101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101111101101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101111101101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10101011111101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10101011110101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101011110101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111111111011110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101111111101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "01111111111001110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "01111111111001110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101111111001110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101111101011110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10101011101111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10101011101101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10111011111101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011111101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011111100110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011111100110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101111101100110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101111101101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101111101101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111111100101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011101101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111111101100110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111111101101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111111101101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111111101101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111111101111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10111111101111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111111101111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111111101111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10111111101111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111111101110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10111011101111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011101111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011101110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011101110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111111101110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10111111101111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10111111101111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10111111101101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10111111101101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10111111101101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10111011111111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011111110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111111101100110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10101111111101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111111111101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111111111100110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111101101100110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101111111101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00101111111101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00101111111101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "01111111111101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "01101111111101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "01111111111001110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "01111111111001110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "01111111111001110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "01111111111101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101011111101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101011111101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011111101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111111111101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011111101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011111100110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011111100110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011111100110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "01111011111100110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101111111110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10101011101111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10111011101101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011101101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011111100110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111111101100110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111111101100110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111111101101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111111100101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111111101101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111111101100110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111111101100110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111111101101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111111101101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111111101101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111111101111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111111101111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10111111101101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111111101111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111111101110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10111111101111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011101110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011101110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10111011111110010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011101110010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10111111101111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10111111101111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111111101100110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111111101101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10111111101101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10111011101111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111111101110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111111101101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111111101101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101111101101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101111101101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101111101101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10101011111101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10101011111101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10111111111101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10111011111101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10111011111101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10111011111101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111111111101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111111111111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "01111011111111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "01111011111110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "01111011111101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101011101101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101111101101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111111101101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111111101100110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101011101101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10101011101101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011111100110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101011111100110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101111111101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101111111101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111111111101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111111101101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111111101100110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101111101101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111111100101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011110101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011100101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111111101100110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011100100110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111111101101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111111101101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111111101101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111111101101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111111100111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10111111101101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111111101101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111111101101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111111101101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011101110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011101110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011101110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111111101110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10111111101111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111111101111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111111101111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111111101101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111111101101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111111101111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111111101100110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111111101101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111111101101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101111101101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101111101101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101111101101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101111101111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101111101111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101101101111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10101111101101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101011101101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10101011101101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10101011111101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10101011111101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10111011111111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10111011111111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10111011111111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101111111101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101111111101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101111111101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101111111001110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101111111111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101111101111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101111101101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101011101101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10101011110101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011111101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011111101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111111111101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111111111100110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111111111101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111111111101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111111110101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111111110101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111111101100110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111111101101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111111101101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111111101101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111111101101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111111101101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10111111101111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111111101101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111111101100110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111111101100110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111111101100110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111111101111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10111111101111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111111111110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111111101110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10111111101101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111111101110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111111101101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10111111101101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10111111111101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011111111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111111101000110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111111101101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111111101101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101111101111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101111101111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101111101111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101111101111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101111101111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101111101111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101111101111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101111100101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101111101101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10101011111101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10101011111101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10111011111101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10101011111101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011111111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "01111111111101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "01111111111101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "01111011111101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "01111011111101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011110101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101111111101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "01101111111101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101111111101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111111111101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111111101101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111111101101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111111101101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101111101101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111111101101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111111100101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011100101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011100101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111111100101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111111101101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111111101101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111111100101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111111100101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111111100101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111111101101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111111101100110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111111101111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111111101111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111111101111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10111111101111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10111111101111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011101110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011101101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011101100110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111111101111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111111101101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10111111101101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10111011101111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011111111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111111111100110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111111101101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10111111111101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111111111101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101111111100110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101111101100110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101111101111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101111101111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101111101111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101111101111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10101111101111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10101111101111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10101011101111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10101011101101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10101011111101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10101011111101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10111011111111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111111111100110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111111111100110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011110101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011110101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011110101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011111101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011111101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011111101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011111101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011111101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "01111011111100110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "01111011111100110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111111111100110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111111111101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101111101101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10111111111111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011111110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011101100110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111111101100110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111111101101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111111101101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111111101101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111111101100110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111111101100110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111111101110010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10111111101111010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111111101111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111111101100010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10111111101111010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10111011101110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10111011101111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10111011101111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10111011111101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011101110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10111111101101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111111101101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10111011101101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011100101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111111100101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111111101111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10111111101101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111111101101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111111101100110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101111101111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101111101101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101111111101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101111111101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101111111101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101111101101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101111101111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101111101111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10101111101111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10101011101111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10101011111101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10111011111111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111111111100110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011111100110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111111110101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101011100101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101111100101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101111101100110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101111101101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101101101101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101111101101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011101101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011101101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011111101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011111100110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111111111100110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101111101101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10111111101101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011111100110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011101100110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111111101101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111111101101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111111101101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111111101100110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111111101100110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111111101100110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10111111101111010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10111011101111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111111101110010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111111101110010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10111011101110010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11011011101110010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10111011101111010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10111011111111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011101110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011101110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10111111100111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10111011101111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011101101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111111101100110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111111101101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10101111111101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00101111111101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10101111111101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011111100110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101111111100110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10101011110101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00101011111101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "01101111111101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "01111111111101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "01111111111100110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "01101111111100110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101111111100110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101111101101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10101011101101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10101011111101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10111011111101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111111111101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101111101100110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101111101100110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101111101101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101111101101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101111101101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101111101101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101111101101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101111101101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101111101101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101111101101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101111101101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111111111101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111111111101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101111101101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10101111101101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10111011111101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011111110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111111101100110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111111101100110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111111101100110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111111101100110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111111101100110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10111111101101010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10111011101101010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011101110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10111011101110010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11011111111110010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11011011101110010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10011011101110010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10111011101111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10111011111111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011101110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111111101110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111111101111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10111011101101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011101100110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111111101100110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111111101101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10101111101101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10111111101101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10111111101101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011101100110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101011101100110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10101111101101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10101011101101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10101011111101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10111011111111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011111101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "01111011111101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "01111011111100110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "01101111111110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101011111101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10101011111101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10101011111101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101111111100110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101111111100110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101111101100110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101111101101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101111100101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101111101101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101111101101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101111101111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101111101101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101111101101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101111101101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10101111101101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101111110101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111111111100110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111111101100110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10101111101101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10111011101101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011101100110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111111101100110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111111101100110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111111101100110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111111101100110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10111111101101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10111011101100110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011111100010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011101110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10011111101111010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11011011111110010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10011111101110010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10111011111110010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11011011101111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10111011101111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011101110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111111101110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10111011101111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10111011111111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111111101100110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111111101101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111111110101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101111110101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101111111101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101111101111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111111101111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101111101111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101111101101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101111101111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101111101111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10101011101101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10101011111101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10111011111101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011111111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "01111011111111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "01111111111100110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "01111011111100110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011111101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101111101100110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101111101100110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101111101101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101111100101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101111100101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101111101111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101111111101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101111111101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101111111101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101111111101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101111101101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101111101111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101111101101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101111101101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111111101101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101111100101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10101111101101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011111100110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011101100110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111111101000110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111111101100110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111111101101010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10111011101101010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10111011101101010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011101100110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111111101110010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10111111111111010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011111110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10111011101111010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10111011101110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11011011101110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011101110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10111111101111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10111111101111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011111110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011101110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111111101110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111111101101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10111111101101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10101011111101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10101011111101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011111101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011111100110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101111110101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10101011111101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00101011111101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "01111111111100110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111111111101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101011111101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10101011111101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10101011111101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10111011111111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111111111111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111111111110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011111110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101111101101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101111111101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "01101111111101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "01111111111101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101111111101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10101111111101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "01111111111101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "01111111111101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "01111111111100110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111111111100110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101111111101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "01101111111101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "01111111111101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111111111100110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111111111100110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101111100101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10101111100101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011111101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011101100110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111111101100110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101111101100110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111111101100110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111111101100010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111111101100110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111111101110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10111111101111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10111011101111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111111101110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10011011101110010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10011011101110010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11011011101110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111111101110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111111100111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10111111101101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011101100110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111111101110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111111101111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111111101101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101111111101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101111101101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111111101111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10101111101101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10111011101101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011101101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10101111101111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10101011111111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10111011111111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "01111011111101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "01111011111100110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011111110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101011111111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10101011111111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10111011111111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10111011111111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111111111101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00101111111101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "01111111111101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111111111100110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111111111100110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101011111100110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10111011111101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10111111111101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111111111101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111111111100110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101111111100110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101111111101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111111111101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111101111100110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111101111100110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111111101110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101111101101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10111111101101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111111101101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011101100110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011101110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111111101101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111111101100110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111111101100110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111111101100110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111111101101010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10101111101111010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011101110010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011101110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10011011101110010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11011011101110010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10011011101111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10111011111111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10111011101111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011101110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111111101100110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111111101110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111111101111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10101111101101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10101011111101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10111011111101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "01111111111100110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111111111110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101111101101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101111111101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101011111101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101011101111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10101011101111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10101011111111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10111011111111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "01111011111111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "01111011111100110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011111110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101011111111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10101011111101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10111011111101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "01111111111101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111111111100110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111101111100110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101111101100110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101011111111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101011101101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101101101101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101101101100110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101101101100110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101111101101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101111101111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101101101110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101101101110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101111101110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101111101111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101111101110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101111101101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101111101101010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10101111101111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011101111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011101100110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111111101100010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111111101101010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111111101100010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10101111101111010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111111101111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011101110010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10011011101110010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11011011101110010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011101111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10111111101111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011111110010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011101110010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011101110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111111101110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111111101111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101011101101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101011111111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10101011101111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10111011111101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10111011111101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011111101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "01101011110110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10101011111101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011111101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011111100110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101011111110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10101011101111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10001011111111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10101011111111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011111111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "01111011111100110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "01111011111100110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011111101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10111011111101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111101111100110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111101111100110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101111111101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "01101111111101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111111111100110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101111111101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101111111101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101111111101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "01111111111001110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "01111111111101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101111111101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101111101101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101111101101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101111101111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101111101111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101111101111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101111101111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101111101111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10101111101111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10111111101111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011101110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10111011101101010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011111111010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011111110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10111111101111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011101110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011101110010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10111011111110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011101110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10111011101111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111111101110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011101110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011101110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011101111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111111101110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111111101111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10101011101111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10101011111101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011111101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011111110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10101011101111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10101011101101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10101011111101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10001011110101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10001011110111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011111111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "01111011111110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011111110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101011111111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10101011111111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10101011111111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011111111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011111110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011111110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011111111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111111111100110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101011111101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101011111100110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101111111100110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101011111101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10101111111101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "01111111111101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111111111101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111111111100110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111111111100110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111111101100110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101111101100110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101111101101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101111101111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101111101111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101111101111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101111101111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111111101111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111111101111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111111101110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111111101111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10111111101101010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011111100110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011111110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011111111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011101110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011101110010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011101110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011101110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011101110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111111101111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111111101111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011101110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101111101110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101111101111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101111101111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101011101111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10101011101111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10101011111101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011111101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "01111011110110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101111111111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10101011111101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10101011110101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10001011110101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10001011110111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10111011111111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "01111011111110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011111110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101011111110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10101011111111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10111011111111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10111011111111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111111111111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011111100110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101011111100110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011111101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011111100110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101111111101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10101111111101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011111101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111111111100110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111101111100110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111111101100110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111111101100110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101111101110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101111101110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101111101111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101111101111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101111101111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111111101111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111111101111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111111101101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111111101101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111111101101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111111101101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10111111101101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111111101101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10111111101111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011101110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111101101110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111111101111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111111101110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111111101110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111111101111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11011111101111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111111101110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10101111101111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10111011101111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111111111111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111111101111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10101011101111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101011111111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101011111111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10111011101101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10111011111101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10101011111111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101011111111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011111110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11001011111101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10001011110111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10001011110111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10111011111111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111111111111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "01111011111110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011111110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101011111111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10111011111111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10111011111111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111111111110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011111101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011111101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011111101010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101111111101010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101111111100110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101101101100110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101111101110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101111101100110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101111101100110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101111101110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101111101111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101111101111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111111101111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101111101111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111111101111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101111101101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101111101101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111111111101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101111101101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101111101100110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111111101100110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111111101101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111111101101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111111101101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111111101110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10111111101111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011101110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011101110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011101110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10111011101111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011111110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11011011101111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101011111110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10111011101111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10011011111111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11011011111110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10101011101111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10101011111111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101011111111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101011111110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10101011101111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10101011101111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10101011110111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011111111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011111110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11001011111111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10001011110111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10001011110111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10011011111111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011111111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011111110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011111110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011111111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10111011111111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011111111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011111101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011111100110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101011111100110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101111101100110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101111101100110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101111101101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101011111101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101111111100110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101111101100110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101111101111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101111101111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111111101011110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101111101111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101111101101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101111101111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101111101111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101111101110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101111101110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101111101110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101111101110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101111101111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111111101111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101111101111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101111101111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111111101111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10111111101111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011101110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10111011101111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011101110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10101011101111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011111110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10101011101111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101011111111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101011101111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10001011111111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11001011111111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011111110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10101011101111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10001011110111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11001011111110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101011111110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10001011111111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10101011101111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10001011110111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011111111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011111110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11001011111111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10001011110111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10101011111111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10111011111111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011111110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011111111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011111110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011111110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10111011111111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111111111100110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101011111100110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101111111100110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101111111100110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101011111101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101111111101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101011111100110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101111101100110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10101111101101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00101111111101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "01111111111101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111111111010110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101111101111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101111101100110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101111101110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101111101110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101111101111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101111101110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101111101111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101111101111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101111101111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101111101111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101111101111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10101111101101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111111101101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10111011111111010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11001011111110010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10101011111111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101011111110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10101011111111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11011011111110010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101011101111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101011111111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101011111110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10101011101111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10101011111111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011111111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11011111111110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10101011101111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101011111111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101011111110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10001011111111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101011111111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10001011110111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10001011110111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011111111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011111110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101011111110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10101011111111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10101011111111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10111011111111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10111111111111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011111110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011111110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011111110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011111100110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "01101011111101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101011111100110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101011111100110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101011111101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101011111101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101011111100110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101011101101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10101111111101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00111011111101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "01111111111100110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111111111100110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101011111100110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101111101100110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101111101111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101111101111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101111101110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101111101111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101111101111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101111101110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101111101110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111111101111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111111101111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111111101101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111111101101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101011111110010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011111111010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10111011111111010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101011111110010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10101011111111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "01011011111110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11001011101111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10011011111111010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11011111111110010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11001011111111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10111011111111010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011111111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011111110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101011111110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10101011101111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011111111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10111011111111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011111110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101011111110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10101011111111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10011011111111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011111110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011111110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011111110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10111011111111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10111011111111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10111011111111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111111111111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011111100110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011111110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00111011111101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011111100110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011111100010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101011111100010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011111100110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "01111011111100110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101011111100010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10101011111101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "01111011111101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011111100110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "01111011111101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011111100110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011111100110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101111101100110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00101011111101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "01101011111100110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101011101100110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101111101111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101111101111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10101111111101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101011111100110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101111101110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10101111101111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10101111111101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101111111100110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101111101100110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10111011101111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011111110010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101011101110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10111011111111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "01011011111110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11001011101111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10011011111111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11011011111110010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11011011111110010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10001011111111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10101011111111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011111110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011111110010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11001011111111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10101011111111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011111110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011111111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011111110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011111111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10101011111111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10111011111111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011111110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011111110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10111011111111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10111011111111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10111011111111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10111011111111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111111111110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111111111111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011111100110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011111100110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101011111100110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011111101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011111101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101011111100010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10111011111101010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10111011111101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011111101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "01111011111101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011111100110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011111100110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011111100110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10101111111101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101011111100110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101011111100110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101111101110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101111111101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101011101110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10101011111101010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101011101100010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101111101111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10101111111111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00111011111111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011111110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101011101110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10101011111111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101011111110010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101011101111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10101011111111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "01011011111110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11011011111110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10111011111111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011111110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11011011111110010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011111110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10101011111111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011111111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11011011111110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11011011110110010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10001011111111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011111111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011111110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10111011111111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011111110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011111110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10111011111111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10111011111111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011111110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011111111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10111011111111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10111011111111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10111011111111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111111111111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10111111111111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10111011111101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10111011111101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011111100110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "01111011111111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011111100110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011111101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10111011111101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011111101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10111011111101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011111100110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011111100110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011111101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00111011111101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "01101011111100110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011111100010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011101100110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10101111111101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011111100110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101011101100110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101111101101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101111101110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10101011101111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10101011111111010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011111110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011111110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101011111111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101011111111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101011111110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101011101111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10001011111111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011111110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011111110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10001011111111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10111011111111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11011011111110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11011011111110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10101011111111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10111011111111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011111110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11011011111110010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10001011111111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10111011111111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011111111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11011011111111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011111111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011111110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10101011111111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10111011111111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011111111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011111110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011111110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10111011111111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10111011111111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10111011111111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10111111111111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10111011111101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111111111100110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10111011111111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011111110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011111100110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011111100110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011111101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10111011111111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011111101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011111100110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011111101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00111011111101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011111110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011111110010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011111110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10101011111101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "01111011111111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011111110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011101110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10101011111111010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101111111110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10101011111111010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10101011111111010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011111110010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011111110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10101011111111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101011111110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101011111110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101011101111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10001011111111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "01111011111111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011111110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10001011111111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10011011111111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011111110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11001011111110010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011111110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10111011111111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011111110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011111110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11011011111110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10001011111111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10111011111111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011111110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10111011111111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011111110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011111110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10111011111111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10111011110111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111111111110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011111110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011111110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10111011111111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10111111111111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10111111111111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111111111100110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111111111111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011111110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011111100110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011111100110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011111100110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011111111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011111111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011111100010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011111101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10111011111101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011111111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011111100110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011111100010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011111111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10101011111101010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011111110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011111110010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10101011111111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "01111011111111010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101011111110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10101011111111010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00011011111111010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011111110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011111110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "01001011111111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11011011111110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101011111110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101011101110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10101011111111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00111011111111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011111110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11011011111111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10111011111111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011111110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11001011111110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011111110010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10111011111111010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10111011111111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011111110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011111110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10011011111111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10111011111111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011111110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011111111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10111011111111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011111110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011111111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10111011111111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10111011111111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011111110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011111110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011111110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10111011111111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10111111111111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111111111100110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111111111100110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011111100110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10111011111101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011111100110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011111110010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10111011111111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011111110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011111101010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10111011111101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "01111011111101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011111110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011111100010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101011111100110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10101011111111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00111011111111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011111110010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011101111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00111011111111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "01111011111110010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101011111111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00111011111111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10111011111110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011111110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011101111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "01101011111111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011111110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011111110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11001011111110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10001011111111010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10011011111111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011111110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11011011111111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10011011111111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11011011111110010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11011011111110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011111110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011111110010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011111111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011111111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11011011111110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10001011111110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10101011111111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011111111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11011011111110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10111011111111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011111110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011111110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10111011111111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10111011111111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10111011111101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011111111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011111110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011111110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10111011111111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011111110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011111100110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10111011111101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10111011111101010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10111011111111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10111011111110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10111011111111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011111110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011111111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10111011111111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111111111110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011111110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10101011111111010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00111011111111010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10111011111111010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011111110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011111110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10111011111111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00111011111111010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11011011111110010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10101011101111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10111011111111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10011011111110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011111110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101011101111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10111011111111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011111110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101011111110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10001011111111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10001011111111010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10011011111111010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011111110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11011011111110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10001011111111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11011011111110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11011011111110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10011011111111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011111110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011111111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10111011111111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011111110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11011011111110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10001011111111010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10111011111111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011111110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011111111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10111011111111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011111110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011111111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10111011111111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10111011111111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10111111111111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111111111110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011111110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011111110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011111110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011111110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10111011111101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10111011111101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10111111111111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10111011111111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011111110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011111110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10111011111111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111111111111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011111110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011111110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00111011111111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10111011111111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10101011111111010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011111110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011111110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10101011111111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011111111010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11011011111110010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10101011111111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10111011111111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011111110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011111110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10111011111111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "01011011111110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11011011111110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11011011111110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10101011111111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10011011111111010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10011011111111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011111110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11011011111110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10011011111111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011111111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011111110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10011011111111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10111011111111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011111110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011111111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011111110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011111110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10101011111111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10111011111111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011111111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011111110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10111011111111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10111011111111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111111111110110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10111011111111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10111011111111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111011111111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111111111101110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111111111111110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11111111111110110000000000000000";
        wait for clk_period;

        new_data <= '0';
        wait for clk_period*10;

        -- #transfers - 1
        new_data <= '1';
        data_input <= "00000000000000000101111010000111";
        wait for clk_period;

        -- Height - 1
        new_data <= '1';
        data_input <= "00000000000000000000000000110110";
        wait for clk_period;

        -- Width - 1
        new_data <= '1';
        data_input <= "00000000000000000000000000110110";
        wait for clk_period;

        -- x_z_slice
        new_data <= '1';
        data_input <= "00000000000000000000011011100000";
        wait for clk_period;

        -- Values
        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '0';
        wait for clk_period*10;

        ----------------------------------
        -- Filters set from DDR to BRAM --
        ----------------------------------
        -- Indices
        -- #filters
        new_data <= '1';
        data_input <= "00000000000000000000000000001000";
        wait for clk_period;

        -- Height - 1
        new_data <= '1';
        data_input <= "00000000000000000000000000000010";
        wait for clk_period;

        -- Width - 1
        new_data <= '1';
        data_input <= "00000000000000000000000000000010";
        wait for clk_period;

        -- Depth
        new_data <= '1';
        data_input <= "00000000000000000000000000100000";
        wait for clk_period;

        -- #transfers
        new_data <= '1';
        data_input <= "00000000000000000000000000001001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00100100101110010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10101100100100010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00100100000010100000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "01001100100100100000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00101111110010000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10000000110010000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00100100000000100000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "01000100000011000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "01001100100001000000000000000000";
        wait for clk_period;

        -- #filters
        new_data <= '1';
        data_input <= "00000000000000000000000000001000";
        wait for clk_period;

        -- Height - 1
        new_data <= '1';
        data_input <= "00000000000000000000000000000010";
        wait for clk_period;

        -- Width - 1
        new_data <= '1';
        data_input <= "00000000000000000000000000000010";
        wait for clk_period;

        -- Depth
        new_data <= '1';
        data_input <= "00000000000000000000000000100000";
        wait for clk_period;

        -- #transfers
        new_data <= '1';
        data_input <= "00000000000000000000000000001001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000100010011010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "01000000011011000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10000100011000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11000000010101000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "01000100001001000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10010001011001000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11010000000001100000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000011000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001010011000000000000000000";
        wait for clk_period;

        -- #filters
        new_data <= '1';
        data_input <= "00000000000000000000000000001000";
        wait for clk_period;

        -- Height - 1
        new_data <= '1';
        data_input <= "00000000000000000000000000000010";
        wait for clk_period;

        -- Width - 1
        new_data <= '1';
        data_input <= "00000000000000000000000000000010";
        wait for clk_period;

        -- Depth
        new_data <= '1';
        data_input <= "00000000000000000000000000100000";
        wait for clk_period;

        -- #transfers
        new_data <= '1';
        data_input <= "00000000000000000000000000001001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10101000101000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10000000000001000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00011010100000010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "01010001000000100000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00101111101100000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000100000100000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00001000110000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001100000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00001000110000000000000000000000";
        wait for clk_period;

        -- #filters
        new_data <= '1';
        data_input <= "00000000000000000000000000001000";
        wait for clk_period;

        -- Height - 1
        new_data <= '1';
        data_input <= "00000000000000000000000000000010";
        wait for clk_period;

        -- Width - 1
        new_data <= '1';
        data_input <= "00000000000000000000000000000010";
        wait for clk_period;

        -- Depth
        new_data <= '1';
        data_input <= "00000000000000000000000000100000";
        wait for clk_period;

        -- #transfers
        new_data <= '1';
        data_input <= "00000000000000000000000000001001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10010100000100000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00101001110100110000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10010101100100000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00010010000110000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "01011111101101100000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00001010100100000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00011011000100000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00001010100100010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10010011000100000000000000000000";
        wait for clk_period;

        -- #filters
        new_data <= '1';
        data_input <= "00000000000000000000000000001000";
        wait for clk_period;

        -- Height - 1
        new_data <= '1';
        data_input <= "00000000000000000000000000000010";
        wait for clk_period;

        -- Width - 1
        new_data <= '1';
        data_input <= "00000000000000000000000000000010";
        wait for clk_period;

        -- Depth
        new_data <= '1';
        data_input <= "00000000000000000000000000100000";
        wait for clk_period;

        -- #transfers
        new_data <= '1';
        data_input <= "00000000000000000000000000001001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00001000110100100000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00101000001010000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00101100101010000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00100000101000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00100000101010100000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00100001000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "01001000000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00001100101000000000000000000000";
        wait for clk_period;

        -- #filters
        new_data <= '1';
        data_input <= "00000000000000000000000000001000";
        wait for clk_period;

        -- Height - 1
        new_data <= '1';
        data_input <= "00000000000000000000000000000010";
        wait for clk_period;

        -- Width - 1
        new_data <= '1';
        data_input <= "00000000000000000000000000000010";
        wait for clk_period;

        -- Depth
        new_data <= '1';
        data_input <= "00000000000000000000000000100000";
        wait for clk_period;

        -- #transfers
        new_data <= '1';
        data_input <= "00000000000000000000000000001001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000001010000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00101010101010000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00100000001010000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10101000101010100000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "01001000100000100000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00001000001000100000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "01100001001100000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00101010100111000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00101000000010100000000000000000";
        wait for clk_period;

        -- #filters
        new_data <= '1';
        data_input <= "00000000000000000000000000001000";
        wait for clk_period;

        -- Height - 1
        new_data <= '1';
        data_input <= "00000000000000000000000000000010";
        wait for clk_period;

        -- Width - 1
        new_data <= '1';
        data_input <= "00000000000000000000000000000010";
        wait for clk_period;

        -- Depth
        new_data <= '1';
        data_input <= "00000000000000000000000000100000";
        wait for clk_period;

        -- #transfers
        new_data <= '1';
        data_input <= "00000000000000000000000000001001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00011010000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000010000100010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00001001000100010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00011010000101000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10010111111000010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "01001010000100010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00011001010100000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00010110010100010000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00011011010000010000000000000000";
        wait for clk_period;

        -- #filters
        new_data <= '1';
        data_input <= "00000000000000000000000000001000";
        wait for clk_period;

        -- Height - 1
        new_data <= '1';
        data_input <= "00000000000000000000000000000010";
        wait for clk_period;

        -- Width - 1
        new_data <= '1';
        data_input <= "00000000000000000000000000000010";
        wait for clk_period;

        -- Depth
        new_data <= '1';
        data_input <= "00000000000000000000000000100000";
        wait for clk_period;

        -- #transfers
        new_data <= '1';
        data_input <= "00000000000000000000000000001001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "10000100000000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00010000000110000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00100001101000000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00101000000010000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "11101010101110100000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00100001000010100000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "01001000001011000000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00101000100010100000000000000000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000000001011100000000000000000";
        wait for clk_period;

        -- Values
        -- #filters
        new_data <= '1';
        data_input <= "00000000000000000000000000001000";
        wait for clk_period;

        -- Height - 1
        new_data <= '1';
        data_input <= "00000000000000000000000000000010";
        wait for clk_period;

        -- Width - 1
        new_data <= '1';
        data_input <= "00000000000000000000000000000010";
        wait for clk_period;

        -- Depth
        new_data <= '1';
        data_input <= "00000000000000000000000000100000";
        wait for clk_period;

        -- #transfers
        new_data <= '1';
        data_input <= "00000000000000000000000000110000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        -- #filters
        new_data <= '1';
        data_input <= "00000000000000000000000000001000";
        wait for clk_period;

        -- Height - 1
        new_data <= '1';
        data_input <= "00000000000000000000000000000010";
        wait for clk_period;

        -- Width - 1
        new_data <= '1';
        data_input <= "00000000000000000000000000000010";
        wait for clk_period;

        -- Depth
        new_data <= '1';
        data_input <= "00000000000000000000000000100000";
        wait for clk_period;

        -- #transfers
        new_data <= '1';
        data_input <= "00000000000000000000000000101000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        -- #filters
        new_data <= '1';
        data_input <= "00000000000000000000000000001000";
        wait for clk_period;

        -- Height - 1
        new_data <= '1';
        data_input <= "00000000000000000000000000000010";
        wait for clk_period;

        -- Width - 1
        new_data <= '1';
        data_input <= "00000000000000000000000000000010";
        wait for clk_period;

        -- Depth
        new_data <= '1';
        data_input <= "00000000000000000000000000100000";
        wait for clk_period;

        -- #transfers
        new_data <= '1';
        data_input <= "00000000000000000000000000100010";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000000";
        wait for clk_period;

        -- #filters
        new_data <= '1';
        data_input <= "00000000000000000000000000001000";
        wait for clk_period;

        -- Height - 1
        new_data <= '1';
        data_input <= "00000000000000000000000000000010";
        wait for clk_period;

        -- Width - 1
        new_data <= '1';
        data_input <= "00000000000000000000000000000010";
        wait for clk_period;

        -- Depth
        new_data <= '1';
        data_input <= "00000000000000000000000000100000";
        wait for clk_period;

        -- #transfers
        new_data <= '1';
        data_input <= "00000000000000000000000000110100";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        -- #filters
        new_data <= '1';
        data_input <= "00000000000000000000000000001000";
        wait for clk_period;

        -- Height - 1
        new_data <= '1';
        data_input <= "00000000000000000000000000000010";
        wait for clk_period;

        -- Width - 1
        new_data <= '1';
        data_input <= "00000000000000000000000000000010";
        wait for clk_period;

        -- Depth
        new_data <= '1';
        data_input <= "00000000000000000000000000100000";
        wait for clk_period;

        -- #transfers
        new_data <= '1';
        data_input <= "00000000000000000000000000011111";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000000";
        wait for clk_period;

        -- #filters
        new_data <= '1';
        data_input <= "00000000000000000000000000001000";
        wait for clk_period;

        -- Height - 1
        new_data <= '1';
        data_input <= "00000000000000000000000000000010";
        wait for clk_period;

        -- Width - 1
        new_data <= '1';
        data_input <= "00000000000000000000000000000010";
        wait for clk_period;

        -- Depth
        new_data <= '1';
        data_input <= "00000000000000000000000000100000";
        wait for clk_period;

        -- #transfers
        new_data <= '1';
        data_input <= "00000000000000000000000000101001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000000000000000000000";
        wait for clk_period;

        -- #filters
        new_data <= '1';
        data_input <= "00000000000000000000000000001000";
        wait for clk_period;

        -- Height - 1
        new_data <= '1';
        data_input <= "00000000000000000000000000000010";
        wait for clk_period;

        -- Width - 1
        new_data <= '1';
        data_input <= "00000000000000000000000000000010";
        wait for clk_period;

        -- Depth
        new_data <= '1';
        data_input <= "00000000000000000000000000100000";
        wait for clk_period;

        -- #transfers
        new_data <= '1';
        data_input <= "00000000000000000000000000101110";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000000000000";
        wait for clk_period;

        -- #filters
        new_data <= '1';
        data_input <= "00000000000000000000000000001000";
        wait for clk_period;

        -- Height - 1
        new_data <= '1';
        data_input <= "00000000000000000000000000000010";
        wait for clk_period;

        -- Width - 1
        new_data <= '1';
        data_input <= "00000000000000000000000000000010";
        wait for clk_period;

        -- Depth
        new_data <= '1';
        data_input <= "00000000000000000000000000100000";
        wait for clk_period;

        -- #transfers
        new_data <= '1';
        data_input <= "00000000000000000000000000101000";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '1';
        data_input <= "00000001000000010000000100000001";
        wait for clk_period;

        new_data <= '0';


        -- while DEBUG_first_done = '0' loop
            -- wait for clk_period;
        -- end loop;
        
        -- report "IDLE";
        -- for i in PUs - 1 downto 0 loop            
            -- write(my_line, to_uint(idle_count(i)));
            -- writeline(output, my_line);
        -- end loop;
        
        -- report "MULT";
        -- for i in PUs - 1 downto 0 loop            
            -- write(my_line, to_uint(mult_count(i)));
            -- writeline(output, my_line);
        -- end loop;
        
        -- assert false report "Simulation finished successfully" severity failure;
 wait;
    end process;
end;